module ALU(ain,bin,sout,zero,overflow,negative);
