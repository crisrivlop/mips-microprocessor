module reg_bank();


endmodule

